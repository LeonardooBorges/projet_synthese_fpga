LIBRARY IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity eInstMem is
	port (
		signal ReadAddr : in std_logic_vector (6 downto 0);
		signal clk : in std_logic;
		signal Instruction31_0 : out std_logic_vector (31 downto 0)
	);
end entity eInstMem;

use work.SpyOnMySigPkg.all;

architecture aInstMem of eInstMem is
type instmem is array (0 TO 31) of std_logic_vector(31 downto 0);
signal mem : instmem := ((("00100000000010000000000011111111"),("10100000000010000000000000000000"),("10000000000010000000000000000000"),("00100000000010010101010000110010"),("00000001000010010100100000100110"),("10101100000010010000000000000000"),("00100000000010110000000000001101"),("00100000000011000000000001000000"),("00000001011011000101100000100101"),("10100000000010110000000000000100"),("00110001011010110000000000000000"),("00100000000010110000000011111001"),("00100000000011000000000000001111"),("00000001011011000101100000100100"),("00110101011010110000000001000000"),("10100000000010110000000000000101"),("00100000000011010100100111111111"),("00000000000011010110101000000010"),("00110101101011010100110100000000"),("00000000000011010110110000000000"),("00110101101011010101000001010011"),("10101100000011010000000000001000"),
others=> (others=>'0'))); --here we put the code that we want to execute





begin
	process (mem)    
	begin
	for i in 0 TO 31 LOOP            
		Globalmem(i) <= mem(i);
	end LOOP;
	end process;

	process (clk)
	begin
	if rising_edge(clk) then
		Instruction31_0 <= mem(to_integer(unsigned(ReadAddr))/4);
	end if;
	end process;
end architecture aInstMem;
